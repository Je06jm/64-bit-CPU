`include "rtl/defines.svh"

//import defines::*;

module MMUTest();

endmodule

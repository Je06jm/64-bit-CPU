`include "rtl/types.svh"
`include "rtl/requests.svh"

module Ld1 #(
    parameter sizeKB = 16
) (
    
);
    
endmodule

`include "rtl/types.svh"
`include "rtl/requests.svh"



`include "rtl/defines.svh"

import defines::*;
